library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity XOR is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end XOR;

architecture rtl of XOR is

begin

end architecture;