-- Write a general sequence detector.